module tb;
reg clk=0,rst;
always begin 
    clk=~clk;
    #50;
    end

Pipeline_top dut(.clk(clk),.rst(rst));
    initial begin 
        $dumpfile("pipeline_top.vcd");
        $dumpvars(0, tb);
    end
    initial begin
        rst<=1'b0;
        #200;
        rst<=1'b1;
        #1000;
    end


    endmodule
